typedef struct packed {
    
}ins_t;