
interface base_iterface();
    // input_1
    // input_2
    // output
endinterface