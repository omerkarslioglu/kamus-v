`include "uvm_macros.svh"

import uvm_pkg::*;

module uvm_tb_top();

    /*
        instantiate our design
    */

    /*
    initial begin
        run_test("our_test");
    end
    */
endmodule